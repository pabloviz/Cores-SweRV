
//General
`define OVI_SBID_WIDTH 5

//Issuing
`define OVI_INSTR_WIDTH 32
`define OVI_SCALAROPND_WIDTH 64
`define OVI_VL_WIDTH 15
`define OVI_SEW_WIDTH 3

//Completing
`define OVI_DATA_WIDTH 64
`define OVI_FFLAGS_WIDTH 5
`define OVI_VSTART_WIDTH 14
