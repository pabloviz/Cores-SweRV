
//General
`define OVI_SBID_WIDTH 5
`define OVI_MEMDATA_WIDTH 512

//Issuing
`define OVI_INSTR_WIDTH 32
`define OVI_SCALAROPND_WIDTH 64
`define OVI_VL_WIDTH 15 //12
`define OVI_SEW_WIDTH 2

//Completing
`define OVI_DATA_WIDTH 64
`define OVI_FFLAGS_WIDTH 5
`define OVI_VSTART_WIDTH 14 //12

//LOAD / STORE packets
`define CPU_PACKET_WIDTH 64 //32 
`define SUBPACKET_BITS ($clog2(`OVI_MEMDATA_WIDTH / `CPU_PACKET_WIDTH)) 
//`define SUBPACKET_BITS_DCCM ($clog2(`OVI_MEMDATA_WIDTH / 32)) 
//`define SUBPACKET_BITS_AXI ($clog2(`OVI_MEMDATA_WIDTH / 64)) 
